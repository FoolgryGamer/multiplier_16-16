module Compressor(
    input ,
    input ,
    input ,
    input ,
    input ,
    output ,
    output ,
    output 
);

endmodule