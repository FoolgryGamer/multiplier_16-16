module multi_top(
    input [15:0] A,
    input [15:0] B,
    output [31:0] out
);




endmodule